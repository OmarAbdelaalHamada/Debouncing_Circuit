module FSM(clk,rst_n,sync_signal,timer_done,debouncer_out,timer_en);
input clk,rst_n,sync_signal,timer_done;
output reg debouncer_out,timer_en;

endmodule