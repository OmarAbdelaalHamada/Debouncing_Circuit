module Debouncing_Circuit();

endmodule